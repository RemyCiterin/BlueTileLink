import Connectable :: *;
import BlockRam :: *;
import TLTypes :: *;
import RegFile :: *;
import Vector :: *;
import Utils :: *;
import AXI4 :: *;
import Fifo :: *;
import Ehr :: *;

`include "TL.defines"

export mkTileLinkClientFSM;

Bool verbose = False;

typedef enum {
  // Ready to receive a new acquire request
  IDLE = 0,

  // Send probe requests, and wait for response
  PROBE_WAIT = 1,

  // Wait for a grant response
  GRANT_WAIT = 2,

  // Receive a probe burst
  PROBE_BURST = 3,

  // Send a grant burst
  GRANT_BURST = 4,

  // Receive a put burst
  PUT_BURST = 5,

  // Send a get burst
  GET_BURST = 6,

  // Receive a release burst
  RELEASE_BURST = 7
} TLClientState deriving(FShow, Eq, Bits);

interface AcquireBuffer#(`TL_ARGS_DECL);
  // Write into the buffer a beat from a cache due to a probe request
  method Action enqProbe(Bit#(dataW) value);

  // Write into the buffer a beat from memory
  method Action enqMem(Bit#(dataW) value);

  // Read one word from the buffer
  method ActionValue#(Bit#(dataW)) deq;

  // Start a new transaction
  method Action start;
endinterface

module mkAcquireBuffer#(Bit#(sizeW) logSize) (AcquireBuffer#(`TL_ARGS));
  Bit#(sizeW) logBusSize = fromInteger(log2(valueOf(dataW)/8));
  Bit#(addrW) maxOffset = (1 << (logSize - logBusSize)) - 1;

  RegFile#(Bit#(addrW), Maybe#(Bit#(dataW))) buffer <- mkRegFile(0, maxOffset);

  function Bit#(addrW) next(Bit#(addrW) idx) = idx == maxOffset ? 0 : idx + 1;
  Reg#(Maybe#(Bit#(addrW))) memHead <- mkReg(Invalid);
  Reg#(Bit#(addrW)) probeHead <- mkReg(0);
  Reg#(Bit#(addrW)) deqHead <- mkReg(0);

  Reg#(Bool) isInit <- mkReg(False);

  rule init if (!isInit);
    buffer.upd(deqHead, Invalid);
    deqHead <= next(deqHead);

    if (deqHead == maxOffset)
      isInit <= True;
  endrule

  method Action enqProbe(Bit#(dataW) value) if (isInit);
    action
      buffer.upd(probeHead, Valid(value));
      probeHead <= next(probeHead);
    endaction
  endmethod

  method Action enqMem(Bit#(dataW) value)
    if (isInit &&& memHead matches tagged Valid .head);
    action
      if (buffer.sub(head) == Invalid && deqHead <= head)
        buffer.upd(head, Valid(value));

      memHead <= head == maxOffset ? Invalid : Valid(head+1);
    endaction
  endmethod

  method ActionValue#(Bit#(dataW)) deq
    if (buffer.sub(deqHead) matches tagged Valid .data);
    buffer.upd(deqHead, Invalid);
    deqHead <= next(deqHead);
    return data;
  endmethod

  method Action start if (memHead == Invalid);
    action
      doAssert(probeHead == 0, "probe head must be 0");
      doAssert(deqHead == 0, "deq head must be 0");
      memHead <= Valid(0);
    endaction
  endmethod
endmodule

// A simple TileLink snoop controller
module mkTileLinkClientFSM#(
    Bit#(sinkW) sink,
    Bit#(sizeW) logSize,
    TLMaster#(`TL_ARGS) master,
    TLSlave#(addrW, dataW, sizeW, sinkW, 0) slave,
    function Bit#(sourceW) repr(Bit#(sourceW) source),
    Vector#(nSource, Bit#(sourceW)) sources
  ) (Empty) provisos (Alias#(Bit#(TAdd#(1, TLog#(nSource))), sourceIdx));

  Reg#(Bool) waitAccessAck <- mkReg(False);

  Bit#(sizeW) logBusSize = fromInteger(log2(valueOf(dataW)/8));

  function Bit#(addrW) align(Bit#(addrW) address);
    return address & ~((1 << logSize) - 1);
  endfunction

  Reg#(TLClientState) state <- mkReg(IDLE);
  Reg#(TLClientState) nextState <- mkReg(IDLE);

  Reg#(ChannelA#(`TL_ARGS)) channelA <- mkReg(?);
  Reg#(TLPerm) acquirePerm <- mkReg(?);

  AcquireBuffer#(`TL_ARGS) buffer <- mkAcquireBuffer(logSize);

  function Action startGrant();
    action
      state <= case (channelA.opcode) matches
        tagged AcquireBlock .* : GRANT_BURST;
        tagged AcquirePerms .* : GRANT_BURST;
        PutData : PUT_BURST;
        GetFull : GET_BURST;
      endcase;
    endaction
  endfunction

  // Release state
  Reg#(TLSize) releaseSize <- mkReg(0);
  Reg#(Bit#(addrW)) releaseAddr <- mkReg(0);

  sourceIdx numSource = fromInteger(valueOf(nSource));

  ProbeFSM#(0, nSource, `TL_ARGS) probeM <- mkProbeFSM(logSize, master, sources);

  // Grant state
  Reg#(Bit#(addrW)) grantSize <- mkReg(0);

  Ehr#(2, Bit#(addrW)) fillAddr <- mkEhr(0);
  Ehr#(2, Bit#(addrW)) fillSize <- mkEhr(0);
  Ehr#(2, Bool) needFill <- mkEhr(False);

  rule receiveChannelA if (state == IDLE && !waitAccessAck);
    let msg = master.channelA.first;

    grantSize <= 1 << logSize;
    master.channelA.deq;
    channelA <= msg;

    if (verbose)
      $display("Client: ", fshow(msg));

    buffer.start();
    fillAddr[0] <= msg.address;
    fillSize[0] <= 1 << logSize;
    needFill[0] <= True;

    doAssert(msg.size == logSize, "Invalid channel A request size");

    Bit#(nSource) srcs = -1;
    for (Integer i=0; i < valueOf(nSource); i = i + 1) begin
      if (sources[i] == repr(msg.source)) srcs[i] = 0;
    end

    if (numSource > 1) begin
      Cap cap = permChannelA(msg.opcode) == T ? N : B;
      probeM.start(?, ProbeBlock(cap), align(msg.address), srcs);
      state <= PROBE_WAIT;
    end else
      state <= GRANT_BURST;
  endrule

  rule probeWrite
    if (
      (state == PROBE_WAIT || state == PROBE_BURST) &&
      (!waitAccessAck || state == PROBE_BURST)
    );

    match {.*, .data, .last} <- probeM.write;

    buffer.enqProbe(data);
    slave.channelA.enq(ChannelA{
      address: channelA.address,
      opcode: PutData,
      data: data,
      size: logSize,
      source: sink,
      mask: -1
    });

    waitAccessAck <= True;

    state <= last ? PROBE_WAIT : PROBE_BURST;
  endrule

  (* preempts = "probeWrite,rresponseMEM" *)
  rule rresponseMEM
    if (
      needFill[0] && fillSize[0] > 0 &&
      slave.channelD.first.source == sink &&
      slave.channelD.first.opcode == AccessAckData
    );
    buffer.enqMem(slave.channelD.first.data);
    slave.channelD.deq;

    fillSize[0] <= fillSize[0] - fromInteger(valueOf(dataW)/8);
    fillAddr[0] <= fillAddr[0] + fromInteger(valueOf(dataW)/8);

    if (fillSize[0] == fromInteger(valueOf(dataW)/8)) begin
      needFill[0] <= False;
    end
  endrule

  rule toGrant if (state == PROBE_WAIT);
    state <= GRANT_BURST;
    probeM.finish;

    slave.channelA.enq(ChannelA{
      address: channelA.address,
      opcode: GetFull,
      size: logSize,
      source: sink,
      mask: ?,
      data: ?
    });
  endrule

  rule sendGrant if (state == GRANT_BURST);
    let data <- buffer.deq;

    Bool last = grantSize == fromInteger(valueOf(dataW)/8);

    master.channelD.enq(ChannelD{
      opcode: GrantData(probeM.exclusive ? T : B),
      source: channelA.source,
      size: channelA.size,
      sink: sink,
      data: data
    });

    if (last) begin
      state <= GRANT_WAIT;
    end

    grantSize <= grantSize - fromInteger(valueOf(dataW)/8);
  endrule

  rule receiveGrantAck
    if (state == GRANT_WAIT && !needFill[1] && master.channelE.first.sink == sink);

    if (verbose)
      $display("Client: ", fshow(master.channelE.first));

    master.channelE.deq;
    state <= IDLE;
  endrule

  rule receiveRelease if (
      (state == IDLE || state == PROBE_WAIT) &&&
      master.channelC.first.opcode matches tagged Release .*
    );

    master.channelC.deq;
    let msg = master.channelC.first;

    doAssert(msg.size == logSize, "Invalid channel C request size");

    master.channelD.enq(ChannelD{
      opcode: ReleaseAck,
      source: msg.source,
      size: msg.size,
      sink: sink,
      data: ?
    });
  endrule

  rule receiveReleaseData if (
      (state == IDLE || state == PROBE_WAIT || state == RELEASE_BURST) &&&
      master.channelC.first.opcode matches tagged ReleaseData .* &&&
      (!waitAccessAck || state == RELEASE_BURST)
    );

    master.channelC.deq;
    let msg = master.channelC.first;
    TLSize size = state == RELEASE_BURST ? releaseSize : 1 << msg.size;
    Bit#(addrW) addr = state == RELEASE_BURST ? releaseAddr : msg.address;
    Bool first = state != RELEASE_BURST;

    doAssert(msg.size == logSize, "Invalid channel C request size");

    if (first) waitAccessAck <= True;
    slave.channelA.enq(ChannelA{
      opcode: PutData,
      data: msg.data,
      address: addr,
      size: logSize,
      source: sink,
      mask: -1
    });

    releaseAddr <= addr + fromInteger(valueOf(dataW)/8);
    releaseSize <= size - fromInteger(valueOf(dataW)/8);
    Bool last = size == fromInteger(valueOf(dataW)/8);

    if (last) begin
      master.channelD.enq(ChannelD{
        opcode: ReleaseAck,
        source: msg.source,
        size: msg.size,
        sink: sink,
        data: ?
      });
    end

    if (first && !last) begin
      state <= RELEASE_BURST;
      nextState <= state;
    end else if (last && !first) begin
      state <= nextState;
    end
  endrule

  rule sendReleaseAck if (
      slave.channelD.first.source == sink &&
      slave.channelD.first.opcode == AccessAck &&
      waitAccessAck
    );

    slave.channelD.deq;
    waitAccessAck <= False;
  endrule
endmodule

// An interface used by a cache to have a TileLink Client interface, can be
// used as example by a Snoop Filter, a LLC, or just a snoop controller
interface ProbeFSM#(numeric type indexW, numeric type nSource, `TL_ARGS_DECL);
  // Request to the FSM to send a probe signal to a set of sources, and write-back the result
  method Action start(Bit#(indexW) idx, OpcodeB op, Bit#(addrW) addr, Bit#(nSource) owners);

  // Write a received data lane to the response buffer
  method ActionValue#(Tuple3#(Bit#(indexW), Bit#(dataW), Bool)) write;

  // Return if any agent still own the data
  method Bool exclusive;

  // Return if we received some data
  method Bool receiveData;

  // Finish th eprobe sequence
  method Action finish;
endinterface

module mkProbeFSM#(
    Bit#(sizeW) logSize,
    TLMaster#(`TL_ARGS) master,
    Vector#(nSource, Bit#(sourceW)) sources
  ) (ProbeFSM#(indexW, nSource, `TL_ARGS))
  provisos (Alias#(Bit#(TAdd#(1, TLog#(nSource))), sourceIdx));

  let metaC <- mkMetaChannelC(master.channelC);
  let channelC = metaC.channel;
  let message = channelC.first;

  sourceIdx numSource = fromInteger(valueOf(nSource));
  Bit#(sizeW) logBusSize = fromInteger(log2(valueOf(dataW)/8));

  Reg#(Bit#(addrW)) address <- mkReg(?);
  Reg#(Bool) exc <- mkReg(True);

  Reg#(Bit#(nSource)) toSend <- mkReg(0);
  Reg#(Bit#(nSource)) toReceive <- mkReg(0);

  Reg#(OpcodeB) opcode <- mkReg(?);
  Reg#(Bit#(indexW)) index <- mkReg(?);
  Reg#(Bool) hasData <- mkReg(?);

  Reg#(Bool) busy <- mkReg(False);

  function sourceIdx findSource(Bit#(sourceW) source);
    sourceIdx idx = ?;

    for (Integer i=0; i < valueOf(nSource); i = i + 1) begin
      if (source == sources[i]) idx = fromInteger(i);
    end

    return idx;
  endfunction

  rule receiveProbeAck
    if (message.opcode matches tagged ProbeAck .reduce);

    let idx = findSource(message.source);
    doAssert(toReceive[idx] == 1, "Receive two ProbeAck from the same source");
    toReceive[idx] <= 0;

    if (verbose)
      $display("Client: ", fshow(message));

    if (reduceTo(reduce) != N) exc <= False;

    channelC.deq;
  endrule

  rule sendProbe if (firstOneFrom(toSend,0) matches tagged Valid .idx);

    let source = sources[idx];
    ChannelB#(`TL_ARGS) msg = ChannelB{
      address: address,
      opcode: opcode,
      source: source,
      size: logSize
    };

    master.channelB.enq(msg);
    toSend[idx] <= 0;
  endrule

  method ActionValue#(Tuple3#(Bit#(indexW), Bit#(dataW), Bool)) write
    if (message.opcode matches tagged ProbeAckData .reduce);

    let idx = findSource(message.source);
    doAssert(toReceive[idx] == 1, "Receive two ProbeAckData from the same source");
    doAssert(!hasData, "Receive a cache block from a Probe request multiple times");
    channelC.deq;

    if (verbose)
      $display("Client: ", fshow(message));

    index <= index + 1;

    if (metaC.last) begin
      if (reduceTo(reduce) != N) exc <= False;
      toReceive[idx] <= 0;
      hasData <= True;
    end

    return tuple3(index, message.data, metaC.last);
  endmethod

  method Action start(Bit#(indexW) idx, OpcodeB op, Bit#(addrW) addr, Bit#(nSource) owners)
    if (!busy);
    action
      exc <= True;
      busy <= True;
      index <= idx;
      opcode <= op;
      address <= addr;
      hasData <= False;
      toSend <= owners;
      toReceive <= owners;
    endaction
  endmethod

  method Action finish if (toReceive == 0 && toSend == 0 && busy);
    action
      busy <= False;
    endaction
  endmethod

  method Bool exclusive = exc;
  method Bool receiveData = hasData;
endmodule
